import axi_pkg::*;
import sauria_pkg::*;
import sauria_addr_pkg::*;
import uvm_pkg::*;

`include "uvm_macros.svh"


