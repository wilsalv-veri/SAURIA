`ifndef SAURIA_SCBD_PKG
`define SAURIA_SCBD_PKG

package sauria_scbd_pkg;

    import uvm_pkg::*;
    import sauria_common_pkg::*;
    import sauria_golden_model_pkg::*;
    
    `include "sauria_dma_req_addr_scbd.sv"

endpackage

`endif //SAURIA_SCBD_PKG