interface sauria_df_controller_ifc;

    logic dma_tile_ptr_advance;
    df_ctrl_substate_t df_ctrl_substate;
    
endinterface