import axi_pkg::*;
import sauria_pkg::*;
import sauria_addr_pkg::*;
import df_ctrl_pkg::*;
import uvm_pkg::*;

`include "uvm_macros.svh"


