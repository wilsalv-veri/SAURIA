class sauria_dma_rd_addr_scbd extends uvm_scoreboard;

    `uvm_component_utils(sauria_dma_rd_addr_scbd)

    string message_id = "SAURIA_DMA_RD_ADDR_SCBD";

    `uvm_analysis_imp_decl(_dma_rd_addr)
    uvm_analysis_imp_dma_rd_addr #(sauria_axi4_rd_addr_seq_item , sauria_dma_rd_addr_scbd) receive_dma_rd_addr;
     
    tensor_ptr_model       ptr_model;
    sauria_computation_params computation_params;

    sauria_axi4_addr_t           tensor_ptr_next_exp_addr;
    sauria_axi4_rd_addr_seq_item dma_rd_addr;

    function new(string name="sauria_dma_rd_addr_scbd", uvm_component parent=null);
        super.new(name,parent);
    endfunction

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        ptr_model       = tensor_ptr_model::type_id::create("tensor_ptr_model");
   
        receive_dma_rd_addr = new("RECEIVE_DMA_RD_ADDR_ANALYSIS_IMP", this);
        
        if (!uvm_config_db #(sauria_computation_params)::get(this, "", "computation_params", computation_params))
            `sauria_info(message_id, "Failed to get access to computation params")
    endfunction

    virtual task run_phase(uvm_phase phase);
        wait_params_to_be_shared();
        ptr_model.configure_model(computation_params);
    endtask

    virtual task wait_params_to_be_shared();
        wait(computation_params.tensors_start_addr_shared);
        wait(computation_params.shared);
    endtask

    function write_dma_rd_addr(sauria_axi4_rd_addr_seq_item dma_rd_addr);
        
        check_model_configured();
        this.dma_rd_addr         = dma_rd_addr;
        tensor_ptr_next_exp_addr = ptr_model.get_next_exp_address();
        check_rd_address();
    endfunction

    virtual function void check_rd_address();
        if(tensor_ptr_next_exp_addr != dma_rd_addr.araddr)
            `sauria_error(message_id, $sformatf("DMA Read Address Mismatch Exp: 0x%0h Act: 0x%0h", tensor_ptr_next_exp_addr, dma_rd_addr.araddr))
    endfunction

    virtual function void check_model_configured();
        if (!(computation_params.tensors_start_addr_shared && computation_params.shared))
            `sauria_fatal(message_id, "Tensor Ptr Model Not Configured Yet. Ignore Results!")
    endfunction

endclass